module ui

pub fn test_input_event_test(){
	a := &InputEvent{}
	println("InputEvent : ${a}")
}
